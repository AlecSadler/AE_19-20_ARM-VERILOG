module msb1 (output [1:3]z,input [1:8]x);

  assign z[1]= x[1] | (!x[1] & x[2]) | (!x[1] & !x[2] & x[3]) | (!x[1] & !x[2] & !x[3] & x[4]);
  assign z[2]= x[1] | (!x[1] & x[2]) | (!x[1] & !x[2] & !x[3] & !x[4] & x[5]) | (!x[1] & !x[2] & !x[3] & !x[4] & !x[5] & x[6]);
  assign z[3]= x[1] | (!x[1] & !x[2] & x[3]) | (!x[1] & !x[2] & !x[3] & !x[4] & x[5]) |
                (!x[1] & !x[2] & !x[3] & !x[4] & !x[5] & !x[6] & x[7]);

endmodule
