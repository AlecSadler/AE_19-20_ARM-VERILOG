module omega (output [0:7]z, input [0:7]s);

  assign z= s;

endmodule
