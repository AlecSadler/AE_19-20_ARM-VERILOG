module omega (output z, input state);

  assign z= state;

endmodule
