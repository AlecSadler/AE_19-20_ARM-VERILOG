module sigma (output [0:7]new_s,input [0:7]s,input x);

  assign new_s[0]= s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x;

  assign new_s[1]= (s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x);

  assign new_s[2]= (s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x);

  assign new_s[3]= (s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x);

  assign new_s[4]= (s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & !s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x);

  assign new_s[5]= (s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & !s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & !s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & s[4] & s[5] & s[6] & s[7] & !x);

  assign new_s[6]= (s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & !s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & !s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & !s[5] & !s[6] & s[7] & x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & s[5] & s[6] & s[7] & !x);

  assign new_s[7]= (s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & !s[2] & s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & !s[5] & s[6] & s[7] & x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & !s[5] & !s[6] & s[7] & x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & s[5] & s[6] & s[7] & !x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & !s[5] & !s[6] & !s[7] & x) |
                   (!s[0] & !s[1] & !s[2] & !s[3] & !s[4] & !s[5] & s[6] & s[7] & !x);

endmodule
